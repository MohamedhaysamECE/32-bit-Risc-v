module adderplus4(
 input [31:0]A,
 output [31:0] Y
 );
 
assign Y = A + 32'd4; 

endmodule
